module calculateStats();

endmodule 